module main

fn main() {
	println(square(3).str())
}

fn square(val int) int {
	return val * val
}
